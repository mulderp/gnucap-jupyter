pulse_ckt.sp
 spice
v1 (1 0) pulse (0 1)

.print tran v(1)
.tran 0 1 .1
.tran trace all

.end
