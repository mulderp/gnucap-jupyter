pulse_ckt.sp
* simple pulse
v1 1 0 pulse iv=0 pv=1 rise=0.3

.print tran v(1)
.tran trace all

.end
