pulse_ckt.sp
* simple pulse
v1 1 0 pulse iv=0 pv=1 delay=0.6 rise=0.1

.print tran v(1)
.tran trace all

.end
