** simulation nmos
Vds 1 0 DC +10V
Vgs 2 0 DC +3V
M1 1 2 0 0 nmos_enhance L=10u W=400u

* model statement (Level 1 by default)
.MODEL nmos_enhance nmos (kp=20u Vto=+2 lambda=0)

** output
.print DC V(1) I(Vds)

** analysis
.DC Vds 0V 3V 100mV
